netcdf empty {
}
